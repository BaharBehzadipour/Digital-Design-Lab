`default_nettype none
`timescale 1ps/1ps
`include "dec4_16.v"

module dec4_16_tb;

reg [3:0] W;
wire [0:15] Y;
reg Enable;

dec4_16 UUT (.W(W),  .Y(Y), .Enable(Enable));

initial begin
    $dumpfile("dec4_16_tb.vcd");
    $dumpvars(0, dec4_16_tb);


    Enable=1;

  if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for En=0");
  #20


    Enable=0;
    W[0] = 0;
    W[1] = 0;
    W[2] = 0;
    W[3] = 0;

            if(Y[0]!=1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 0000");
  #20

  Enable=0;
    W[0] = 1;
    W[1] = 0;
    W[2] = 0;
    W[3] = 0;

  if(Y[0]==1 || Y[1]!=1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 0001");
  #20

    Enable=0;
    W[0] = 0;
    W[1] = 1;
    W[2] = 0;
    W[3] = 0;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]!=1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 0010");
  #20

    Enable=0;
    W[0] = 1;
    W[1] = 1;
    W[2] = 0;
    W[3] = 0;

            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]!=1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 0011");
  #20

    Enable=0;
    W[0] = 0;
    W[1] = 0;
    W[2] = 1;
    W[3] = 0;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]!=1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 0100");
  #20


    Enable=0;
    W[0] = 1;
    W[1] = 0;
    W[2] = 1;
    W[3] = 0;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]!=1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 0101");
  #20

    Enable=0;
    W[0] = 0;
    W[1] = 1;
    W[2] = 1;
    W[3] = 0;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]!=1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 0110");
  #20

    Enable=0;
    W[0] = 1;
    W[1] = 1;
    W[2] = 1;
    W[3] = 0;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]!=1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 0111");
  #20

    Enable=0;
    W[0] = 0;
    W[1] = 0;
    W[2] = 0;
    W[3] = 1;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]!=1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 1000");
  #20  


      Enable=0;
    W[0] = 1;
    W[1] = 0;
    W[2] = 0;
    W[3] = 1;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]!=1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 1001");
  #20  


        Enable=0;
    W[0] = 0;
    W[1] = 1;
    W[2] = 0;
    W[3] = 1;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]!=1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 1010");
  #20  

    Enable=0;
    W[0] = 1;
    W[1] = 1;
    W[2] = 0;
    W[3] = 1;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]!=1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 1011");
  #20  

      Enable=0;
    W[0] = 0;
    W[1] = 0;
    W[2] = 1;
    W[3] = 1;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]!=1 ||Y[13]==1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 1100");
  #20  


    Enable=0;
    W[0] = 1;
    W[1] = 0;
    W[2] = 1;
    W[3] = 1;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]!=1 ||Y[14]==1 ||Y[15]==1)
    $display("test fail for 1101");
  #20  

      Enable=0;
    W[0] = 0;
    W[1] = 1;
    W[2] = 1;
    W[3] = 1;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]!=1 ||Y[15]==1)
    $display("test fail for 1110");
  #20  


      Enable=0;
    W[0] = 1;
    W[1] = 1;
    W[2] = 1;
    W[3] = 1;
 
            if(Y[0]==1 || Y[1]==1 || Y[2]==1 ||Y[3]==1 ||Y[4]==1 ||Y[5]==1 ||Y[6]==1 ||Y[7]==1 ||Y[8]==1 ||
  Y[9]==1 ||Y[10]==1 ||Y[11]==1 ||Y[12]==1 ||Y[13]==1 ||Y[14]==1 ||Y[15]!=1)
    $display("test fail for 1111");
  #20  

    $display("*******complete*******");
   
end

endmodule
